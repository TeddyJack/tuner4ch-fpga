// для своевременного вычитывания пакетов из буферов, необходимо, чтобы F_read >= (4 x F_write_max), а лучше (5 x F_write_max)

`include "defines.v"

module source_switch(		// здесь сформировать give_me_one_packet для каждого источника
input SYS_CLK,
input RST,
input [3:0] GOT_FULL_PACKET,

input [31:0] DATA_IN_BUS,

input [7:0] SPI_ADDRESS,
input [7:0] SPI_DATA,
input RISING_SS,

output reg [3:0] RD_REQ,

output reg [7:0] DATA_OUT,
output DCLK_OUT,
output reg D_VALID_OUT,
output reg P_SYNC_OUT

);

//reg [7:0] header_3d_array [3:0][3:0];		// 
//reg [7:0] src;										// число, номер источника
//initial
//begin
//for(src=0; src<4; src=src+1'b1)
//	begin
//	header_3d_array[src][0] = src;			// PLP ID
//	header_3d_array[src][1] = src + 8'd2;	// stream source
//	header_3d_array[src][2] = 8'h00;			// reserved
//	header_3d_array[src][3] = 8'h00;			// reserved
//	end
//end
reg [7:0] header_2d_array [15:0];		// 
reg [7:0] src;										// число, номер источника
initial
begin
for(src=0; src<4; src=src+1'b1)
	begin
	header_2d_array[(src<<2) + 2'h0] = src;			// PLP ID				// (<<2) = (*4)
	header_2d_array[(src<<2) + 2'h1] = src + 8'd2;	// stream source
	header_2d_array[(src<<2) + 2'h2] = 8'h00;			// reserved
	header_2d_array[(src<<2) + 2'h3] = 8'h00;			// reserved
	end
end



assign DCLK_OUT = SYS_CLK;
wire [7:0] DATA_IN [3:0];

genvar i;
generate
for(i=0; i<4; i=i+1)
	begin: wow
	assign DATA_IN[i] = DATA_IN_BUS[(8*i+7):(8*i)];
	end
endgenerate

reg [1:0] state;
parameter [1:0] check_source		= 2'h0;
parameter [1:0] fill_header		= 2'h1;
parameter [1:0] forward_packet	= 2'h2;

reg [1:0] source_counter;
reg [7:0] byte_counter;

always@(posedge SYS_CLK or negedge RST)
begin
if(!RST)
	begin
	source_counter <= 0;
	state <= check_source;
	byte_counter <= 0;
	DATA_OUT <= 0;
	P_SYNC_OUT <= 0;
	RD_REQ <= 4'b0000;
	D_VALID_OUT <= 0;
	end
else
	case(state)
	check_source:
		begin
		D_VALID_OUT <= 0;
		if(GOT_FULL_PACKET[source_counter])
			begin
			state <= fill_header;
			end
		else
			source_counter <= source_counter + 1'b1;
		end
	fill_header:
		begin
		DATA_OUT <= header_2d_array[(source_counter<<2) + byte_counter];	// (<<2) = (*4)
		if(byte_counter < 4)
			begin
			byte_counter <= byte_counter + 1'b1;
			D_VALID_OUT <= 1;
			end
		else
			begin
			byte_counter <= 0;
			D_VALID_OUT <= 0;
			state <= forward_packet;
			end
		end
	forward_packet:
		begin
		D_VALID_OUT <= RD_REQ[source_counter];
		DATA_OUT <= DATA_IN[source_counter];
		if(byte_counter < 8'd188)
			begin
			
			RD_REQ[source_counter] <= 1;
			byte_counter <= byte_counter + 1'b1;
			if(byte_counter == 8'd0)
				P_SYNC_OUT <= 1;
			else
				P_SYNC_OUT <= 0;
			end
		else
			begin
			byte_counter <= 0;
			RD_REQ[source_counter] <= 0;
			source_counter <= source_counter + 1'b1;
			state <= check_source;
			end
		end
	endcase
end

always@(posedge SYS_CLK)
begin
if(RISING_SS && (SPI_ADDRESS >= `ADDR_HEADR_FIRST) && (SPI_ADDRESS <= `ADDR_HEADR_LAST))
	header_2d_array[SPI_ADDRESS-`ADDR_HEADR_FIRST] <= SPI_DATA;
end


endmodule
